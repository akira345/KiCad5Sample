.title KiCad schematic
Q1 GND Net-_D1-Pad1_ Net-_Q1-Pad3_ 2SC1815
R2 +5V Net-_D1-Pad2_ 100
R1 Net-_Q1-Pad3_ Net-_R1-Pad2_ 7.5k
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ LED
SW1 +5V Net-_R1-Pad2_ SW_Push
J1 +5V GND Conn_01x02_Male
.end
